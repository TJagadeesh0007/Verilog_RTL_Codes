module xor_gate(input a,b, output y);

	xor g1(y,a,b);   //Pimitive Gate
	
	//assign y = a^b;
	
endmodule
	
